library verilog;
use verilog.vl_types.all;
entity Tester is
end Tester;
